module adder8 (); 

endmodule
